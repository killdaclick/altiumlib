***************** Power Discrete MOSFET Electrical Parameters ***********************
** Product: FQD12N20L
** Package: D-PAK
**-----------------------------------------------------------------------------------
.SUBCKT FQD12N20L 20 10 30
Rg  10 1 1.58
M1  2 1 3 3 DMOS L=1u W=1u
.MODEL DMOS NMOS (VTO={1.84*{-0.00096*TEMP+1.024}} KP={TEMP*0.0072+15.6}
+ THETA=0.08  VMAX=4.0E5  LEVEL=3) 
Cgs 1 3 813p
Rd  20 4 0.092  TC=0.009
Dds 3 4 DDS
.MODEL DDS D(BV={200*{0.000875*TEMP+0.978125}} M=0.52 CJO=1260p VJ=0.58)
Dbody 3 20 DBODY
.MODEL DBODY  D(IS=1.8E-12  N=1.0  RS=0.0079  EG=1.06  TT=154n)
Ra  4 2  0.092 TC=0.009
Rs  3 5  0.011
Ls  5 30 1.97n
M2  1 8 6 6 INTER
E2  8 6 4 1 2
.MODEL INTER NMOS(VTO=0  KP=10  LEVEL=1)
Cgdmax 7 4 630p
Rcgd 7 4 10meg
Dgd  6 4 DGD
Rdgd 4 6 10meg
.MODEL DGD D(M=0.42  CJO=630p  VJ=0.18)
M3  7  9 1 1 INTER
E3  9  1 4 1 -2
.ENDS

********************* Power Discrete MOSFET Thermal Model **********************
.SUBCKT FQD12N20L_Thermal TH TL
CTHERM1 TH 6 1.20e-5
CTHERM2 6 5  3.10e-4
CTHERM3 5 4  3.00e-3
CTHERM4 4 3  3.40e-2
CTHERM5 3 2  1.70e-1
CTHERM6 2 TL 1.80e-1 
RTHERM1 TH 6 8.20e-3
RTHERM2 6 5  1.80e-2
RTHERM3 5 4  3.04e-1
RTHERM4 4 3  4.50e-1
RTHERM5 3 2  6.50e-1
RTHERM6 2 TL 8.40e-1
.ENDS FQD12N20L_Thermal 
**-----------------------------------------------------------------------------------
** Creation: Oct.-31-2007
** Fairchild Semiconductor

