.SUBCKT MSS1278-105 1 2
R2 1 3 1.7
RVAR1 3 4 {8.10E-03}
LVAR 4 2 {1000uH}
C1 3 5 13.20pF
R1 5 2 90
.ENDS
