*DEVICE=BZX84C6V2,D

* BZX84C6V2 D model
* created using Parts release 7.1 on 03/30/98 at 14:50
* Parts is a MicroSim product.
.MODEL BZX84C6V2 D
+ IS=110.88E-18
+ N=.92657
+ RS=.85899
+ IKF=149.75
+ CJO=108.46E-12
+ M=.34501
+ VJ=.72044
+ ISR=48.986E-9
+ BV=6.3329
+ IBV=1.0062
+ TT=121.76E-9
*$
