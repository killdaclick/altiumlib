*==============================================
*P-EMOS 3T pinout: D,G,S
*Copyright (c) 1996 MicroCode Engineering, Inc.
*All Rights Reserved
*
*See other copyright notices at end of file.
*==============================================

*PMOS
*Default P-Channel MOSFET parameter values
.MODEL MPMOS~ PMOS()

*IRF9640  MCE  4-2-96
*200V  11A  .5 ohms HEXFET pkg:TO-220 2,1,3
.SUBCKT XIRF9640  10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  .236
RS  30  3  13.5M
RG  20  2  16.3
CGS  2  3  1.11N
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  1.04N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 THETA=60M VMAX=416K ETA=2M VTO=-3 KP=2.46)
.MODEL DCGD D (CJO=1.04N VJ=.6 M=.68)
.MODEL DSUB D (IS=45.6N N=1.5 RS=.386 BV=200 CJO=1.24N VJ=.8 M=.42 TT=250N)
.MODEL DLIM D (IS=100U)
.ENDS XIRF9640


*   Copyright notice for all models labeled "ZETEX":
*
*                          (C)  1992 ZETEX PLC
*
*   The copyright in these models  and  the designs embodied belong
*   to Zetex PLC ("Zetex").  They  are  supplied  free of charge by
*   Zetex for the purpose of research and design and may be used or
*   copied intact  (including this notice)  for  that purpose only.
*   All other rights are reserved. The models are believed accurate
*   but  no condition  or warranty  as to their  merchantability or
*   fitness for purpose is given and no liability in respect of any
*   use is accepted by Zetex PLC, its distributors or agents.
*
*
*   Zetex PLC, Fields New Road, Chadderton, Oldham  OL9 8NP  U.K.
