*FQD7P20 200V P-CHANNEL DMOSFET ELECTRICAL PARAMETERS

*------------------------------------------------------------------------------------

.SUBCKT  FQD7P20   20  10  30

Rg     10    1    1

M1      2    1    3    3    DMOS    L=1u   W=1u

.MODEL DMOS PMOS (VTO={-3.9 * (-0.00088*TEMP+1.022)} KP={4.4 * (-0.00012*TEMP+1.003)}

+ THETA=0.04    VMAX=1.52E5   LEVEL=3)

Cgs 1   3   680P

Rd  20  4   236m   TC=0.00083

Dds 4   3   DDS

.MODEL DDS D(BV={200*(0.0008*TEMP+0.98)}  M=0.5      CJO=115p   VJ=0.8)

Dbody   20  3   DBODY

.MODEL DBODY D(IS=1.2E-13    N=1.05     RS=96.3m    EG=1.17    TT=180n)

Ra 4    2   110m   TC=0.00083

Rs 3    5   11m    

Ls 5    30  1.0n

M2 1    8   6    6   INTER

E2 8    6   4    1   2

.MODEL INTER PMOS (VTO=0   KP=10   LEVEL=1)

Cgdmax  7  4    925P

Rcgd    7  4    10meg

Dgd     4  6    DGD

Rdgd    4  6    10meg

.MODEL DGD D(M=0.74   CJO=925P    VJ=0.62)

M3      7  9  1  1  INTER

E3      9  1  4  1  -2

.ENDS FQD7P20

*-------------------------------------------------------------------------------------

*FAIRCHILD      CASE: D-PAK      PID: FQD7P20 

*NOV-18-2000 CREATION  

