**************** Power Discrete MOSFET Electrical Circuit Model *****************
** Product Name: 2N7002
** Package: TO-236AB
** 60V N-Channel MOSFET
**-------------------------------------------------------------------------------
.SUBCKT F2N7002  20  10  30
Rg 10  1  1.58
M1 2   1  3   3  DMOS   L=1u  W=1u
.MODEL DMOS NMOS (VTO={2.10*{-0.00064*TEMP+1.016}}  KP={{-0.0319*TEMP}+1.022}
+ THETA=0.04  VMAX=5.0E5  ETA=0.001  LEVEL=3)
Cgs   1   3    16p
Rd    20  4    0.13  TC=0.0067
Dds   3   4    DDS
.MODEL  DDS  D(BV={60*{0.000775*TEMP+0.980625}}  M=0.38  CJO=25p  VJ=0.48)
Dbody 3   20    DBODY
.MODEL DBODY  D(IS=3.0E-14  N=1.0  RS=2.015  EG=1.16  TT=52n)
Ra    4    2    0.13 TC=0.0067
Rs    3    5    0.01
Ls    5    30   1.0n
M2    1    8    6    6   INTER
E2    8    6    4    1   2
.MODEL INTER  NMOS(VTO=0  KP=10  LEVEL=1)
Cgdmax 7   4    46p
Rcgd   7   4    10meg
Dgd    6   4    DGD
Rdgd   4   6    10meg
.MODEL DGD D(M=0.56  CJO=46p  VJ=0.384)
M3     7   9   1    1   INTER
E3     9   1   4    1   -2
.ENDS

**-------------------------------------------------------------------------------
** Creation: Nov.-05-2007   Rev: 0.0
** Fairchild Semiconductor

